library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.types_encoder.all;
use work.utils_encoder.all;

-- Package Declaration Section
package comp_encoder is

end package comp_encoder;