--------------------------------------------------------------------------------
-- University:	NTNU Trondheim
-- Project:		CCSDS123 Issue 2
-- Engineer:	Cristian Gil Morales
-- Date:		25/02/2021
--------------------------------------------------------------------------------
-- IP name:		metadata_encod
--
-- Description: Defines the "Encoder Metadata" from compressed image header part
--
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package metadata_encod is


end package metadata_encod;