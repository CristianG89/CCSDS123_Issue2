library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.types.all;
use work.utils.all;

-- Package Declaration Section
package comp_encoder is

end package comp_encoder;