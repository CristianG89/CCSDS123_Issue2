library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.types_image.all;

-- Package Declaration Section
package hybrid_code_table is	
	
	type hybrid_code_table_t is record
		-- input_code	: array_unsigned_t;
		output_code	: array_integer_t;
		output_size	: array_integer_t;
	end record hybrid_code_table_t;
	
	subtype hybrid_code_table0_t is hybrid_code_table_t (
		-- input_code(104 downto 0),
		output_code(104 downto 0),
		output_size(104 downto 0)
	);
	
	constant hybrid_code_table0_c : hybrid_code_table0_t := (
		-- input_code  => (x"00", x"010", x"011", x"012", x"013", x"014", x"015", x"016", x"017", x"018", x"019", x"01A", x"01B", x"01C", x"01X", x"020", x"021", x"022", x"023", x"024", x"025", x"026", x"027", x"028", x"029", x"02A", x"02B", x"02C", x"02X", x"03", x"04", x"05", x"06", x"07", x"08", x"09", x"0A", x"0B", x"0C", x"0X", x"1", x"2", x"3", x"40", x"41", x"42", x"43", x"440", x"441", x"442", x"443", x"444", x"445", x"446", x"447", x"448", x"449", x"44A", x"44B", x"44C", x"44X", x"45", x"46", x"47", x"48", x"49", x"4A", x"4B", x"4C", x"4X", x"5", x"6", x"70", x"71", x"72", x"73", x"74", x"75", x"76", x"77", x"78", x"79", x"7A", x"7B", x"7C", x"7X", x"80", x"81", x"82", x"83", x"84", x"85", x"86", x"87", x"88", x"89", x"8A", x"8B", x"8C", x"8X", x"9", x"A", x"B", x"C", x"X"),
		output_code => (16#19#, 16#57#, 16#d7#, 16#37#, 16#af#, 16#1af#, 16#6f#, 16#16f#, 16#3f#, 16#23f#, 16#17f#, 16#57f#, 16#1ff#, 16#9ff#, 16#37f#, 16#b7#, 16#77#, 16#f7#, 16#ef#, 16#1ef#, 16#1f#, 16#11f#, 16#13f#, 16#33f#, 16#77f#, 16#ff#, 16#5ff#, 16#dff#, 16#4ff#, 16#15#, 16#35#, 16#d#, 16#2d#, 16#13#, 16#53#, 16#3b#, 16#bb#, 16#f#, 16#10f#, 16#7b#, 16#0#, 16#4#, 16#2#, 16#1d#, 16#3d#, 16#3#, 16#23#, 16#9f#, 16#19f#, 16#5f#, 16#bf#, 16#2bf#, 16#1bf#, 16#3bf#, 16#2ff#, 16#6ff#, 16#3ff#, 16#bff#, 16#fff#, 16#1fff#, 16#7ff#, 16#33#, 16#73#, 16#fb#, 16#7#, 16#8f#, 16#18f#, 16#4f#, 16#14f#, 16#87#, 16#6#, 16#e#, 16#b#, 16#4b#, 16#2b#, 16#47#, 16#c7#, 16#27#, 16#a7#, 16#cf#, 16#1cf#, 16#15f#, 16#35f#, 16#7f#, 16#47f#, 16#df#, 16#6b#, 16#1b#, 16#5b#, 16#67#, 16#e7#, 16#17#, 16#97#, 16#2f#, 16#12f#, 16#2df#, 16#1df#, 16#27f#, 16#67f#, 16#3df#, 16#1#, 16#11#, 16#5#, 16#25#, 16#9#),
		output_size => (5, 8, 8, 8, 9, 9, 9, 9, 10, 10, 11, 11, 12, 12, 11, 8, 8, 8, 9, 9, 9, 9, 10, 10, 11, 11, 12, 12, 11, 6, 6, 6, 6, 7, 7, 8, 8, 9, 9, 8, 3, 3, 3, 6, 6, 6, 6, 9, 9, 9, 10, 10, 10, 10, 11, 11, 12, 12, 13, 13, 12, 7, 7, 8, 8, 9, 9, 9, 9, 8, 4, 4, 7, 7, 7, 8, 8, 8, 8, 9, 9, 10, 10, 11, 11, 10, 7, 7, 7, 8, 8, 8, 8, 9, 9, 10, 10, 11, 11, 10, 5, 5, 6, 6, 5)
	);
	
	subtype hybrid_code_table1_t is hybrid_code_table_t (
		-- input_code(143 downto 0),
		output_code(143 downto 0),
		output_size(143 downto 0)
	);
	
	constant hybrid_code_table1_c : hybrid_code_table1_t := (
		-- input_code  => (x"000", x"001", x"002", x"003", x"004", x"005", x"006", x"007", x"008", x"009", x"00A", x"00X", x"01", x"02", x"030", x"031", x"032", x"033", x"034", x"035", x"036", x"037", x"038", x"039", x"03A", x"03X", x"040", x"041", x"042", x"043", x"044", x"045", x"046", x"047", x"048", x"049", x"04A", x"04X", x"05", x"06", x"07", x"08", x"09", x"0A", x"0X", x"10", x"11", x"12", x"130", x"131", x"132", x"133", x"134", x"135", x"136", x"137", x"138", x"139", x"13A", x"13X", x"14", x"150", x"151", x"152", x"153", x"154", x"155", x"156", x"157", x"158", x"159", x"15A", x"15X", x"160", x"161", x"162", x"163", x"164", x"165", x"166", x"167", x"168", x"169", x"16A", x"16X", x"17", x"18", x"19", x"1A", x"1X", x"20", x"21", x"22", x"230", x"231", x"232", x"233", x"234", x"235", x"236", x"237", x"238", x"239", x"23A", x"23X", x"24", x"250", x"251", x"252", x"253", x"254", x"255", x"256", x"257", x"258", x"259", x"25A", x"25X", x"26", x"27", x"28", x"29", x"2A", x"2X", x"3", x"4", x"5", x"6", x"7", x"8", x"9", x"A0", x"A1", x"A2", x"A3", x"A4", x"A5", x"A6", x"A7", x"A8", x"A9", x"AA", x"AX", x"X"),
		output_code => (16#73#, 16#b#, 16#4b#, 16#9b#, 16#5b#, 16#137#, 16#b7#, 16#11f#, 16#31f#, 16#63f#, 16#13f#, 16#53f#, 16#e#, 16#1e#, 16#db#, 16#3b#, 16#bb#, 16#1b7#, 16#77#, 16#177#, 16#f7#, 16#9f#, 16#33f#, 16#57f#, 16#d7f#, 16#73f#, 16#7b#, 16#fb#, 16#7#, 16#1f7#, 16#f#, 16#10f#, 16#29f#, 16#bf#, 16#4bf#, 16#37f#, 16#b7f#, 16#2bf#, 16#1d#, 16#3d#, 16#13#, 16#53#, 16#e7#, 16#1e7#, 16#2b#, 16#1#, 16#11#, 16#9#, 16#87#, 16#47#, 16#c7#, 16#8f#, 16#18f#, 16#19f#, 16#39f#, 16#6bf#, 16#1bf#, 16#77f#, 16#f7f#, 16#ff#, 16#3#, 16#4f#, 16#14f#, 16#cf#, 16#5f#, 16#25f#, 16#15f#, 16#5bf#, 16#8ff#, 16#4ff#, 16#3ff#, 16#13ff#, 16#cff#, 16#1cf#, 16#2f#, 16#12f#, 16#35f#, 16#df#, 16#3bf#, 16#7bf#, 16#2ff#, 16#aff#, 16#bff#, 16#1bff#, 16#7ff#, 16#ab#, 16#6b#, 16#17#, 16#117#, 16#97#, 16#19#, 16#5#, 16#15#, 16#27#, 16#a7#, 16#67#, 16#af#, 16#1af#, 16#2df#, 16#1df#, 16#7f#, 16#47f#, 16#6ff#, 16#eff#, 16#1ff#, 16#23#, 16#6f#, 16#16f#, 16#ef#, 16#3df#, 16#3f#, 16#27f#, 16#67f#, 16#9ff#, 16#5ff#, 16#17ff#, 16#fff#, 16#1fff#, 16#33#, 16#eb#, 16#1b#, 16#197#, 16#57#, 16#157#, 16#0#, 16#4#, 16#2#, 16#a#, 16#6#, 16#16#, 16#d#, 16#d7#, 16#1d7#, 16#37#, 16#1ef#, 16#3ef#, 16#1f#, 16#21f#, 16#23f#, 16#17f#, 16#dff#, 16#1dff#, 16#97f#, 16#2d#),
		output_size => (7, 7, 7, 8, 8, 9, 9, 10, 10, 11, 11, 11, 5, 5, 8, 8, 8, 9, 9, 9, 9, 10, 11, 12, 12, 11, 8, 8, 8, 9, 9, 9, 10, 11, 11, 12, 12, 11, 6, 6, 7, 7, 9, 9, 8, 5, 5, 5, 8, 8, 8, 9, 9, 10, 10, 11, 11, 12, 12, 12, 6, 9, 9, 9, 10, 10, 10, 11, 12, 12, 13, 13, 12, 9, 9, 9, 10, 10, 11, 11, 12, 12, 13, 13, 13, 8, 8, 9, 9, 9, 5, 5, 5, 8, 8, 8, 9, 9, 10, 10, 11, 11, 12, 12, 12, 6, 9, 9, 9, 10, 10, 11, 11, 12, 12, 13, 13, 13, 7, 8, 8, 9, 9, 9, 3, 3, 4, 4, 5, 5, 6, 9, 9, 9, 10, 10, 10, 10, 11, 12, 13, 13, 12, 6)
	);
	
	subtype hybrid_code_table2_t is hybrid_code_table_t (
		-- input_code(117 downto 0),
		output_code(117 downto 0),
		output_size(117 downto 0)
	);
	
	constant hybrid_code_table2_c : hybrid_code_table2_t := (
		-- input_code  => (x"0", x"10", x"110", x"111", x"112", x"113", x"114", x"115", x"116", x"117", x"118", x"11X", x"120", x"121", x"122", x"123", x"124", x"125", x"126", x"127", x"128", x"12X", x"130", x"131", x"132", x"133", x"134", x"135", x"136", x"137", x"138", x"13X", x"140", x"141", x"142", x"143", x"144", x"145", x"146", x"147", x"148", x"14X", x"15", x"16", x"17", x"18", x"1X", x"200", x"201", x"202", x"203", x"204", x"205", x"206", x"207", x"208", x"20X", x"210", x"211", x"212", x"213", x"214", x"215", x"216", x"217", x"218", x"21X", x"22", x"230", x"231", x"232", x"233", x"234", x"235", x"236", x"237", x"238", x"23X", x"240", x"241", x"242", x"243", x"244", x"245", x"246", x"247", x"248", x"24X", x"25", x"26", x"27", x"28", x"2X", x"3", x"4", x"50", x"51", x"52", x"53", x"54", x"55", x"56", x"57", x"58", x"5X", x"60", x"61", x"62", x"63", x"64", x"65", x"66", x"67", x"68", x"6X", x"7", x"8", x"X"),
		output_code => (16#0#, 16#1#, 16#7d#, 16#3#, 16#43#, 16#3b#, 16#bb#, 16#cf#, 16#1cf#, 16#3bf#, 16#7bf#, 16#7f#, 16#23#, 16#63#, 16#13#, 16#7b#, 16#fb#, 16#2f#, 16#12f#, 16#47f#, 16#27f#, 16#67f#, 16#53#, 16#7#, 16#87#, 16#af#, 16#1af#, 16#df#, 16#2df#, 16#2ff#, 16#aff#, 16#6ff#, 16#47#, 16#c7#, 16#27#, 16#6f#, 16#16f#, 16#1df#, 16#3df#, 16#eff#, 16#1ff#, 16#9ff#, 16#35#, 16#75#, 16#6b#, 16#f7#, 16#1f7#, 16#15#, 16#33#, 16#73#, 16#a7#, 16#67#, 16#ef#, 16#1ef#, 16#17f#, 16#57f#, 16#37f#, 16#b#, 16#4b#, 16#2b#, 16#e7#, 16#17#, 16#1f#, 16#11f#, 16#77f#, 16#ff#, 16#4ff#, 16#9#, 16#97#, 16#57#, 16#d7#, 16#9f#, 16#19f#, 16#3f#, 16#23f#, 16#5ff#, 16#dff#, 16#3ff#, 16#37#, 16#b7#, 16#77#, 16#5f#, 16#15f#, 16#13f#, 16#33f#, 16#bff#, 16#7ff#, 16#fff#, 16#d#, 16#4d#, 16#eb#, 16#f#, 16#10f#, 16#2#, 16#6#, 16#25#, 16#2d#, 16#6d#, 16#1b#, 16#9b#, 16#8f#, 16#18f#, 16#bf#, 16#4bf#, 16#2bf#, 16#1d#, 16#5d#, 16#3d#, 16#5b#, 16#db#, 16#4f#, 16#14f#, 16#6bf#, 16#1bf#, 16#5bf#, 16#19#, 16#39#, 16#5#),
		output_size => (2, 4, 7, 7, 7, 8, 8, 9, 9, 11, 11, 11, 7, 7, 7, 8, 8, 9, 9, 11, 11, 11, 7, 8, 8, 9, 9, 10, 10, 12, 12, 12, 8, 8, 8, 9, 9, 10, 10, 12, 12, 12, 7, 7, 8, 9, 9, 6, 7, 7, 8, 8, 9, 9, 11, 11, 11, 7, 7, 7, 8, 8, 9, 9, 11, 11, 11, 5, 8, 8, 8, 9, 9, 10, 10, 12, 12, 12, 8, 8, 8, 9, 9, 10, 10, 12, 12, 12, 7, 7, 8, 9, 9, 3, 3, 6, 7, 7, 8, 8, 9, 9, 11, 11, 11, 7, 7, 7, 8, 8, 9, 9, 11, 11, 11, 6, 6, 6)
	);
	
	subtype hybrid_code_table3_t is hybrid_code_table_t (
		-- input_code(119 downto 0),
		output_code(119 downto 0),
		output_size(119 downto 0)
	);
	
	constant hybrid_code_table3_c : hybrid_code_table3_t := (
		-- input_code  => (x"000", x"0010", x"0011", x"0012", x"0013", x"0014", x"0015", x"0016", x"001X", x"0020", x"0021", x"0022", x"0023", x"0024", x"0025", x"0026", x"002X", x"003", x"004", x"005", x"006", x"00X", x"01", x"02", x"03", x"04", x"05", x"06", x"0X", x"1", x"20", x"210", x"2110", x"2111", x"2112", x"2113", x"2114", x"2115", x"2116", x"211X", x"212", x"213", x"214", x"215", x"216", x"21X", x"220", x"2210", x"2211", x"2212", x"2213", x"2214", x"2215", x"2216", x"221X", x"222", x"223", x"224", x"225", x"226", x"22X", x"230", x"231", x"232", x"233", x"234", x"235", x"236", x"23X", x"24", x"25", x"26", x"2X", x"30", x"310", x"311", x"312", x"313", x"314", x"315", x"316", x"31X", x"320", x"321", x"322", x"323", x"324", x"325", x"326", x"32X", x"33", x"34", x"35", x"36", x"3X", x"40", x"410", x"411", x"412", x"413", x"414", x"415", x"416", x"41X", x"42", x"43", x"44", x"45", x"46", x"4X", x"5", x"60", x"61", x"62", x"63", x"64", x"65", x"66", x"6X", x"X"),
		output_code => (16#19#, 16#4b#, 16#17#, 16#97#, 16#ef#, 16#1ef#, 16#37f#, 16#77f#, 16#9ff#, 16#2b#, 16#57#, 16#d7#, 16#1f#, 16#11f#, 16#ff#, 16#4ff#, 16#5ff#, 16#43#, 16#23#, 16#18f#, 16#4f#, 16#14f#, 16#2#, 16#a#, 16#1e#, 16#1#, 16#2d#, 16#6d#, 16#6b#, 16#0#, 16#6#, 16#35#, 16#37#, 16#9f#, 16#19f#, 16#23f#, 16#13f#, 16#dff#, 16#3ff#, 16#fff#, 16#63#, 16#3b#, 16#bb#, 16#2df#, 16#1df#, 16#1bf#, 16#d#, 16#b7#, 16#5f#, 16#15f#, 16#33f#, 16#bf#, 16#bff#, 16#7ff#, 16#1fff#, 16#13#, 16#7b#, 16#fb#, 16#3df#, 16#3f#, 16#5bf#, 16#53#, 16#7#, 16#87#, 16#cf#, 16#1cf#, 16#3bf#, 16#7bf#, 16#aff#, 16#25#, 16#eb#, 16#1b#, 16#9b#, 16#11#, 16#33#, 16#47#, 16#c7#, 16#2f#, 16#12f#, 16#7f#, 16#47f#, 16#6ff#, 16#73#, 16#27#, 16#a7#, 16#af#, 16#1af#, 16#27f#, 16#67f#, 16#eff#, 16#1d#, 16#5d#, 16#77#, 16#177#, 16#f7#, 16#9#, 16#b#, 16#67#, 16#e7#, 16#6f#, 16#16f#, 16#17f#, 16#57f#, 16#1ff#, 16#15#, 16#3d#, 16#7d#, 16#1f7#, 16#f#, 16#df#, 16#e#, 16#3#, 16#5b#, 16#db#, 16#10f#, 16#8f#, 16#2bf#, 16#6bf#, 16#2ff#, 16#5#),
		output_size => (5, 7, 8, 8, 9, 9, 11, 11, 12, 7, 8, 8, 9, 9, 11, 11, 12, 7, 7, 9, 9, 9, 4, 4, 5, 5, 7, 7, 8, 2, 4, 6, 8, 9, 9, 10, 10, 12, 12, 13, 7, 8, 8, 10, 10, 11, 6, 8, 9, 9, 10, 10, 12, 12, 13, 7, 8, 8, 10, 10, 11, 7, 8, 8, 9, 9, 11, 11, 12, 6, 8, 8, 8, 5, 7, 8, 8, 9, 9, 11, 11, 12, 7, 8, 8, 9, 9, 11, 11, 12, 7, 7, 9, 9, 9, 5, 7, 8, 8, 9, 9, 11, 11, 12, 6, 7, 7, 9, 9, 10, 5, 7, 8, 8, 9, 9, 11, 11, 12, 6)
	);
	
	subtype hybrid_code_table4_t is hybrid_code_table_t (
		-- input_code(91 downto 0),
		output_code(91 downto 0),
		output_size(91 downto 0)
	);
	
	constant hybrid_code_table4_c : hybrid_code_table4_t := (
		-- input_code  => (x"000", x"0010", x"0011", x"0012", x"0013", x"0014", x"0015", x"0016", x"001X", x"002", x"003", x"004", x"005", x"006", x"00X", x"0100", x"0101", x"0102", x"0103", x"0104", x"0105", x"0106", x"010X", x"0110", x"0111", x"0112", x"0113", x"0114", x"0115", x"0116", x"011X", x"0120", x"0121", x"0122", x"0123", x"0124", x"0125", x"0126", x"012X", x"013", x"014", x"015", x"016", x"01X", x"020", x"0210", x"0211", x"0212", x"0213", x"0214", x"0215", x"0216", x"021X", x"0220", x"0221", x"0222", x"0223", x"0224", x"0225", x"0226", x"022X", x"023", x"024", x"025", x"026", x"02X", x"030", x"031", x"032", x"033", x"034", x"035", x"036", x"03X", x"040", x"041", x"042", x"043", x"044", x"045", x"046", x"04X", x"05", x"06", x"0X", x"1", x"2", x"3", x"4", x"5", x"6", x"X"),
		output_code => (16#5#, 16#3#, 16#2b#, 16#6b#, 16#11f#, 16#9f#, 16#8ff#, 16#4ff#, 16#cff#, 16#d#, 16#33#, 16#73#, 16#1ef#, 16#15f#, 16#35f#, 16#23#, 16#1b#, 16#5b#, 16#19f#, 16#5f#, 16#2ff#, 16#aff#, 16#6ff#, 16#3b#, 16#f7#, 16#f#, 16#13f#, 16#33f#, 16#eff#, 16#1dff#, 16#3ff#, 16#7b#, 16#8f#, 16#4f#, 16#bf#, 16#2bf#, 16#1ff#, 16#13ff#, 16#bff#, 16#e7#, 16#17#, 16#df#, 16#2df#, 16#17f#, 16#1d#, 16#7#, 16#cf#, 16#2f#, 16#1bf#, 16#3bf#, 16#9ff#, 16#1bff#, 16#7ff#, 16#47#, 16#af#, 16#6f#, 16#7f#, 16#27f#, 16#17ff#, 16#fff#, 16#1fff#, 16#97#, 16#57#, 16#1df#, 16#57f#, 16#37f#, 16#b#, 16#d7#, 16#37#, 16#1f#, 16#3df#, 16#77f#, 16#f7f#, 16#5ff#, 16#4b#, 16#b7#, 16#77#, 16#3f#, 16#23f#, 16#ff#, 16#15ff#, 16#dff#, 16#a7#, 16#67#, 16#ef#, 16#0#, 16#2#, 16#1#, 16#9#, 16#13#, 16#53#, 16#27#),
		output_size => (4, 6, 7, 7, 9, 9, 12, 12, 12, 5, 7, 7, 9, 10, 10, 6, 7, 7, 9, 9, 12, 12, 12, 7, 8, 8, 10, 10, 12, 13, 13, 7, 8, 8, 10, 10, 12, 13, 13, 8, 8, 10, 10, 11, 5, 7, 8, 8, 10, 10, 12, 13, 13, 7, 8, 8, 10, 10, 13, 13, 13, 8, 8, 10, 11, 11, 7, 8, 8, 9, 10, 12, 12, 13, 7, 8, 8, 10, 10, 12, 13, 13, 8, 8, 9, 2, 2, 4, 4, 7, 7, 8)
	);
	
	subtype hybrid_code_table5_t is hybrid_code_table_t (
		-- input_code(115 downto 0),
		output_code(115 downto 0),
		output_size(115 downto 0)
	);
	
	constant hybrid_code_table5_c : hybrid_code_table5_t := (
		-- input_code  => (x"0", x"1", x"2000", x"200100", x"200101", x"200102", x"200103", x"200104", x"20010X", x"20011", x"20012", x"20013", x"20014", x"2001X", x"20020", x"20021", x"20022", x"20023", x"20024", x"2002X", x"2003", x"2004", x"200X", x"201000", x"201001", x"201002", x"201003", x"201004", x"20100X", x"20101", x"20102", x"20103", x"20104", x"2010X", x"2011", x"2012", x"2013", x"2014", x"201X", x"20200", x"20201", x"20202", x"20203", x"20204", x"2020X", x"2021", x"2022", x"2023", x"2024", x"202X", x"203", x"204", x"20X", x"210000", x"210001", x"210002", x"210003", x"210004", x"21000X", x"21001", x"21002", x"21003", x"21004", x"2100X", x"2101", x"2102", x"2103", x"2104", x"210X", x"2110", x"2111", x"2112", x"2113", x"2114", x"211X", x"2120", x"2121", x"2122", x"2123", x"2124", x"212X", x"213", x"214", x"21X", x"22000", x"22001", x"22002", x"22003", x"22004", x"2200X", x"2201", x"2202", x"2203", x"2204", x"220X", x"2210", x"2211", x"2212", x"2213", x"2214", x"221X", x"222", x"223", x"224", x"22X", x"23", x"240", x"241", x"242", x"243", x"244", x"24X", x"2X", x"3", x"4", x"X"),
		output_code => (16#0#, 16#1#, 16#b#, 16#1f#, 16#1df#, 16#3df#, 16#5ff#, 16#15ff#, 16#1fff#, 16#4f#, 16#14f#, 16#d7f#, 16#37f#, 16#7ff#, 16#57#, 16#cf#, 16#1cf#, 16#b7f#, 16#77f#, 16#27ff#, 16#177#, 16#2df#, 16#4bf#, 16#11f#, 16#3f#, 16#23f#, 16#dff#, 16#1dff#, 16#3fff#, 16#2f#, 16#12f#, 16#f7f#, 16#ff#, 16#17ff#, 16#fb#, 16#7#, 16#2bf#, 16#6bf#, 16#1ff#, 16#d7#, 16#af#, 16#1af#, 16#8ff#, 16#4ff#, 16#37ff#, 16#87#, 16#47#, 16#1bf#, 16#5bf#, 16#11ff#, 16#7b#, 16#1b7#, 16#19f#, 16#9f#, 16#13f#, 16#33f#, 16#3ff#, 16#13ff#, 16#7fff#, 16#6f#, 16#16f#, 16#cff#, 16#2ff#, 16#fff#, 16#c7#, 16#27#, 16#3bf#, 16#7bf#, 16#9ff#, 16#a7#, 16#f7#, 16#1f7#, 16#a7f#, 16#67f#, 16#2bff#, 16#67#, 16#f#, 16#10f#, 16#e7f#, 16#17f#, 16#1bff#, 16#39f#, 16#5f#, 16#bf#, 16#37#, 16#ef#, 16#1ef#, 16#aff#, 16#6ff#, 16#2fff#, 16#e7#, 16#17#, 16#7f#, 16#47f#, 16#19ff#, 16#97#, 16#8f#, 16#18f#, 16#97f#, 16#57f#, 16#3bff#, 16#3b#, 16#25f#, 16#15f#, 16#27f#, 16#5b#, 16#77#, 16#35f#, 16#df#, 16#eff#, 16#1eff#, 16#bff#, 16#b7#, 16#3#, 16#13#, 16#1b#),
		output_size => (1, 2, 5, 9, 10, 10, 13, 13, 14, 9, 9, 12, 12, 14, 8, 9, 9, 12, 12, 14, 9, 10, 11, 9, 10, 10, 13, 13, 15, 9, 9, 12, 12, 14, 8, 8, 11, 11, 13, 8, 9, 9, 12, 12, 14, 8, 8, 11, 11, 13, 8, 9, 10, 9, 10, 10, 13, 13, 15, 9, 9, 12, 12, 14, 8, 8, 11, 11, 13, 8, 9, 9, 12, 12, 14, 8, 9, 9, 12, 12, 14, 10, 10, 11, 8, 9, 9, 12, 12, 14, 8, 8, 11, 11, 13, 8, 9, 9, 12, 12, 14, 7, 10, 10, 12, 7, 9, 10, 10, 13, 13, 14, 9, 5, 5, 7)
	);

	subtype hybrid_code_table6_t is hybrid_code_table_t (
		-- input_code(100 downto 0),
		output_code(100 downto 0),
		output_size(100 downto 0)
	);
	
	constant hybrid_code_table6_c : hybrid_code_table6_t := (
		-- input_code  => (x"0000", x"000100", x"000101", x"000102", x"000103", x"000104", x"00010X", x"00011", x"00012", x"00013", x"00014", x"0001X", x"000200", x"000201", x"000202", x"000203", x"000204", x"00020X", x"00021", x"00022", x"00023", x"00024", x"0002X", x"0003", x"0004", x"000X", x"00100", x"00101", x"00102", x"00103", x"00104", x"0010X", x"0011", x"0012", x"0013", x"0014", x"001X", x"002", x"003", x"004", x"00X", x"01", x"020", x"0210", x"0211", x"0212", x"0213", x"0214", x"021X", x"022", x"023", x"024", x"02X", x"03", x"04", x"0X", x"10", x"1100", x"1101", x"1102", x"1103", x"1104", x"110X", x"111", x"112", x"113", x"114", x"11X", x"12", x"13", x"14", x"1X", x"200", x"20100", x"20101", x"20102", x"20103", x"20104", x"2010X", x"2011", x"2012", x"2013", x"2014", x"201X", x"202", x"203", x"204", x"20X", x"21", x"22", x"23", x"24", x"2X", x"30", x"31", x"32", x"33", x"34", x"3X", x"4", x"X"),
		output_code => (16#2#, 16#13#, 16#4f#, 16#cf#, 16#6ff#, 16#eff#, 16#2fff#, 16#3b#, 16#7b#, 16#47f#, 16#27f#, 16#3ff#, 16#33#, 16#2f#, 16#af#, 16#1ff#, 16#9ff#, 16#1fff#, 16#7#, 16#47#, 16#67f#, 16#aff#, 16#13ff#, 16#5f#, 16#15f#, 16#7bf#, 16#15#, 16#27#, 16#67#, 16#17f#, 16#57f#, 16#bff#, 16#1d#, 16#3d#, 16#2bf#, 16#7f#, 16#1dff#, 16#6#, 16#57#, 16#d7#, 16#3f#, 16#0#, 16#e#, 16#3#, 16#37#, 16#b7#, 16#f7f#, 16#ff#, 16#17ff#, 16#d#, 16#23f#, 16#13f#, 16#37f#, 16#4b#, 16#2b#, 16#16f#, 16#4#, 16#23#, 16#77#, 16#f7#, 16#8ff#, 16#4ff#, 16#37ff#, 16#1b#, 16#5b#, 16#3bf#, 16#b7f#, 16#dff#, 16#9#, 16#ef#, 16#1ef#, 16#1bf#, 16#1#, 16#17#, 16#df#, 16#1df#, 16#1bff#, 16#7ff#, 16#7fff#, 16#f#, 16#8f#, 16#cff#, 16#2ff#, 16#fff#, 16#2d#, 16#33f#, 16#bf#, 16#77f#, 16#19#, 16#5#, 16#1f#, 16#11f#, 16#5bf#, 16#6b#, 16#9f#, 16#19f#, 16#5ff#, 16#15ff#, 16#3fff#, 16#b#, 16#6f#),
		output_size => (3, 6, 8, 8, 12, 12, 14, 7, 7, 11, 11, 13, 6, 8, 8, 12, 12, 14, 7, 7, 11, 12, 13, 9, 9, 11, 5, 7, 7, 11, 11, 13, 6, 6, 10, 11, 13, 4, 8, 8, 10, 3, 4, 6, 8, 8, 12, 12, 14, 6, 10, 10, 12, 7, 7, 9, 3, 6, 8, 8, 12, 12, 14, 7, 7, 11, 12, 13, 5, 9, 9, 11, 4, 7, 9, 9, 13, 13, 15, 8, 8, 12, 12, 14, 6, 10, 10, 12, 5, 5, 9, 9, 11, 7, 9, 9, 13, 13, 15, 7, 9)
	);

	subtype hybrid_code_table7_t is hybrid_code_table_t (
		-- input_code(80 downto 0),
		output_code(80 downto 0),
		output_size(80 downto 0)
	);
	
	constant hybrid_code_table7_c : hybrid_code_table7_t := (
		-- input_code  => (x"00", x"0100", x"01010", x"01011", x"01012", x"01013", x"01014", x"0101X", x"01020", x"01021", x"01022", x"01023", x"01024", x"0102X", x"0103", x"0104", x"010X", x"011", x"012", x"013", x"014", x"01X", x"020", x"021", x"0220", x"0221", x"0222", x"0223", x"0224", x"022X", x"023", x"024", x"02X", x"03", x"04", x"0X", x"1000", x"10010", x"10011", x"10012", x"10013", x"10014", x"1001X", x"10020", x"10021", x"10022", x"10023", x"10024", x"1002X", x"1003", x"1004", x"100X", x"101", x"102", x"103", x"104", x"10X", x"110", x"111", x"1120", x"1121", x"1122", x"1123", x"1124", x"112X", x"113", x"114", x"11X", x"12", x"13", x"14", x"1X", x"2", x"30", x"31", x"32", x"33", x"34", x"3X", x"4", x"X"),
		output_code => (16#0#, 16#d#, 16#77#, 16#15f#, 16#df#, 16#17ff#, 16#57ff#, 16#7fff#, 16#f#, 16#1df#, 16#3bf#, 16#37ff#, 16#77ff#, 16#17fff#, 16#1ff#, 16#9ff#, 16#3bff#, 16#2b#, 16#1b#, 16#4ff#, 16#cff#, 16#13ff#, 16#5#, 16#3b#, 16#37#, 16#9f#, 16#19f#, 16#27ff#, 16#67ff#, 16#5fff#, 16#2ff#, 16#aff#, 16#33ff#, 16#1ef#, 16#1f#, 16#27f#, 16#3#, 16#4f#, 16#3f#, 16#13f#, 16#fff#, 16#4fff#, 16#3fff#, 16#2f#, 16#bf#, 16#7f#, 16#2fff#, 16#6fff#, 16#ffff#, 16#5ff#, 16#dff#, 16#7ff#, 16#7#, 16#27#, 16#6ff#, 16#eff#, 16#bff#, 16#17#, 16#6f#, 16#5f#, 16#77f#, 16#ff#, 16#dfff#, 16#1bfff#, 16#3ffff#, 16#2bff#, 16#1bff#, 16#9fff#, 16#b#, 16#67f#, 16#17f#, 16#3ff#, 16#1#, 16#11f#, 16#57f#, 16#37f#, 16#1fff#, 16#bfff#, 16#1ffff#, 16#ef#, 16#1bf#),
		output_size => (1, 4, 7, 9, 9, 15, 15, 17, 7, 9, 10, 15, 15, 17, 12, 12, 14, 6, 6, 12, 12, 14, 4, 6, 7, 9, 9, 15, 15, 16, 12, 12, 14, 9, 9, 11, 4, 7, 9, 9, 15, 15, 16, 7, 9, 10, 15, 15, 17, 12, 12, 14, 6, 6, 12, 12, 14, 6, 8, 9, 11, 11, 16, 17, 18, 14, 14, 16, 6, 11, 11, 13, 3, 9, 11, 11, 16, 17, 18, 9, 10)
	);

	subtype hybrid_code_table8_t is hybrid_code_table_t (
		-- input_code(87 downto 0),
		output_code(87 downto 0),
		output_size(87 downto 0)
	);
	
	constant hybrid_code_table8_c : hybrid_code_table8_t := (
		-- input_code  => (x"0000000000", x"0000000001", x"000000000200", x"000000000201", x"000000000202", x"00000000020X", x"00000000021", x"00000000022", x"0000000002X", x"000000000X", x"000000001", x"000000002", x"00000000X", x"0000000100", x"0000000101", x"0000000102", x"000000010X", x"000000011", x"000000012", x"00000001X", x"000000020", x"000000021", x"000000022", x"00000002X", x"0000000X", x"0000001", x"000000200", x"000000201", x"000000202", x"00000020X", x"00000021", x"00000022", x"0000002X", x"000000X", x"000001", x"000002", x"00000X", x"000010", x"000011", x"000012", x"00001X", x"000020", x"000021", x"000022", x"00002X", x"0000X", x"0001", x"000200", x"000201", x"000202", x"00020X", x"000210", x"000211", x"000212", x"00021X", x"00022", x"0002X", x"000X", x"001", x"002", x"00X", x"010", x"011", x"012", x"01X", x"02", x"0X", x"100", x"101", x"102", x"10X", x"110", x"111", x"112", x"11X", x"12", x"1X", x"200", x"201", x"202", x"20X", x"210", x"211", x"212", x"21X", x"22", x"2X", x"X"),
		output_code => (16#0#, 16#b#, 16#37#, 16#27f#, 16#17f#, 16#3fff#, 16#3bf#, 16#7f#, 16#5fff#, 16#dff#, 16#3#, 16#23#, 16#6ff#, 16#2b#, 16#df#, 16#1df#, 16#1fff#, 16#1f#, 16#11f#, 16#37ff#, 16#13#, 16#9f#, 16#19f#, 16#6fff#, 16#2ff#, 16#1d#, 16#33#, 16#5f#, 16#15f#, 16#fff#, 16#ef#, 16#1ef#, 16#17ff#, 16#4ff#, 16#9#, 16#19#, 16#37f#, 16#5#, 16#f7#, 16#f#, 16#1bff#, 16#15#, 16#8f#, 16#4f#, 16#7ff#, 16#1bf#, 16#1#, 16#d#, 16#cf#, 16#2f#, 16#27ff#, 16#af#, 16#77f#, 16#ff#, 16#ffff#, 16#77#, 16#bff#, 16#2bf#, 16#c#, 16#2#, 16#3f#, 16#a#, 16#3b#, 16#7b#, 16#3ff#, 16#4#, 16#16f#, 16#6#, 16#7#, 16#47#, 16#5ff#, 16#27#, 16#23f#, 16#13f#, 16#2fff#, 16#1b#, 16#1ff#, 16#e#, 16#67#, 16#17#, 16#13ff#, 16#57#, 16#33f#, 16#bf#, 16#7fff#, 16#5b#, 16#9ff#, 16#6f#),
		output_size => (3, 6, 7, 10, 10, 15, 10, 10, 15, 12, 6, 6, 11, 6, 9, 9, 15, 9, 9, 14, 6, 9, 9, 15, 11, 5, 6, 9, 9, 14, 9, 9, 14, 11, 5, 5, 11, 5, 8, 8, 13, 5, 8, 8, 14, 10, 4, 5, 8, 8, 14, 8, 11, 11, 16, 8, 13, 10, 4, 4, 10, 4, 7, 7, 13, 4, 9, 4, 7, 7, 12, 7, 10, 10, 15, 7, 12, 4, 7, 7, 13, 7, 10, 10, 16, 7, 12, 9)
	);

	subtype hybrid_code_table9_t is hybrid_code_table_t (
		-- input_code(105 downto 0),
		output_code(105 downto 0),
		output_size(105 downto 0)
	);
	
	constant hybrid_code_table9_c : hybrid_code_table9_t := (
		-- input_code  => (x"00000000000", x"000000000010", x"000000000011", x"000000000012", x"00000000001X", x"00000000002", x"0000000000X", x"000000000100", x"000000000101", x"000000000102", x"00000000010X", x"00000000011", x"00000000012", x"0000000001X", x"0000000002", x"000000000X", x"000000001000", x"000000001001", x"000000001002", x"00000000100X", x"00000000101", x"00000000102", x"0000000010X", x"0000000011", x"0000000012", x"000000001X", x"0000000020", x"0000000021", x"0000000022", x"000000002X", x"00000000X", x"00000001", x"0000000200", x"0000000201", x"0000000202", x"000000020X", x"000000021", x"000000022", x"00000002X", x"0000000X", x"0000001", x"0000002000", x"0000002001", x"0000002002", x"000000200X", x"000000201", x"000000202", x"00000020X", x"00000021", x"00000022", x"0000002X", x"000000X", x"000001", x"000002", x"00000X", x"000010", x"000011", x"000012", x"00001X", x"00002", x"0000X", x"000100", x"000101", x"000102", x"00010X", x"00011", x"00012", x"0001X", x"00020", x"00021", x"00022", x"0002X", x"000X", x"001000", x"001001", x"001002", x"00100X", x"00101", x"00102", x"0010X", x"0011", x"0012", x"001X", x"00200", x"00201", x"00202", x"0020X", x"0021", x"0022", x"002X", x"00X", x"01", x"02000", x"02001", x"02002", x"0200X", x"0201", x"0202", x"020X", x"021", x"022", x"02X", x"0X", x"1", x"2", x"X"),
		output_code => (16#0#, 16#3b#, 16#1bf#, 16#3bf#, 16#17fff#, 16#1b#, 16#bff#, 16#7#, 16#7f#, 16#27f#, 16#ffff#, 16#33f#, 16#bf#, 16#3fff#, 16#13#, 16#3ff#, 16#27#, 16#17f#, 16#37f#, 16#1ffff#, 16#19f#, 16#2bf#, 16#bfff#, 16#9f#, 16#df#, 16#9fff#, 16#33#, 16#2df#, 16#1df#, 16#7fff#, 16#dff#, 16#3#, 16#b#, 16#3df#, 16#3f#, 16#5fff#, 16#1f#, 16#15f#, 16#efff#, 16#5ff#, 16#1d#, 16#2b#, 16#23f#, 16#13f#, 16#dfff#, 16#11f#, 16#35f#, 16#1fff#, 16#1ef#, 16#25f#, 16#6fff#, 16#9ff#, 16#9#, 16#19#, 16#1ff#, 16#5#, 16#12f#, 16#af#, 16#77ff#, 16#e#, 16#6ff#, 16#15#, 16#1af#, 16#6f#, 16#fff#, 16#b7#, 16#10f#, 16#17ff#, 16#1e#, 16#8f#, 16#18f#, 16#2fff#, 16#2ff#, 16#d#, 16#16f#, 16#ef#, 16#4fff#, 16#77#, 16#4f#, 16#57ff#, 16#97#, 16#57#, 16#47ff#, 16#1#, 16#14f#, 16#cf#, 16#afff#, 16#d7#, 16#1f7#, 16#27ff#, 16#4ff#, 16#6#, 16#11#, 16#1cf#, 16#2f#, 16#37ff#, 16#37#, 16#f#, 16#67ff#, 16#17#, 16#f7#, 16#7ff#, 16#ff#, 16#2#, 16#a#, 16#5f#),
		output_size => (2, 6, 10, 10, 17, 6, 12, 6, 10, 10, 17, 10, 10, 16, 6, 12, 6, 10, 10, 17, 9, 10, 16, 9, 10, 16, 6, 10, 10, 17, 12, 5, 6, 10, 10, 16, 9, 10, 16, 12, 5, 6, 10, 10, 16, 9, 10, 16, 9, 10, 16, 12, 5, 5, 12, 5, 9, 9, 15, 5, 11, 5, 9, 9, 15, 8, 9, 15, 5, 9, 9, 16, 11, 5, 9, 9, 15, 8, 9, 15, 8, 8, 15, 5, 9, 9, 16, 8, 9, 15, 11, 4, 5, 9, 9, 15, 8, 9, 15, 8, 9, 15, 11, 4, 4, 10)
	);

	subtype hybrid_code_table10_t is hybrid_code_table_t (
		-- input_code(102 downto 0),
		output_code(102 downto 0),
		output_size(102 downto 0)
	);
	
	constant hybrid_code_table10_c : hybrid_code_table10_t := (
		-- input_code  => (x"000000000", x"000000001000", x"000000001001", x"000000001002", x"00000000100X", x"00000000101", x"00000000102", x"0000000010X", x"0000000011", x"0000000012", x"000000001X", x"0000000020", x"0000000021", x"0000000022", x"000000002X", x"00000000X", x"000000010000", x"000000010001", x"000000010002", x"00000001000X", x"00000001001", x"00000001002", x"0000000100X", x"0000000101", x"0000000102", x"000000010X", x"000000011", x"000000012", x"00000001X", x"0000000200", x"0000000201", x"0000000202", x"000000020X", x"000000021", x"000000022", x"00000002X", x"0000000X", x"0000001", x"000000200", x"000000201", x"000000202", x"00000020X", x"00000021", x"00000022", x"0000002X", x"000000X", x"000001", x"000002000", x"000002001", x"000002002", x"00000200X", x"00000201", x"00000202", x"0000020X", x"0000021", x"0000022", x"000002X", x"00000X", x"00001", x"000020000", x"000020001", x"000020002", x"00002000X", x"00002001", x"00002002", x"0000200X", x"0000201", x"0000202", x"000020X", x"000021", x"000022", x"00002X", x"0000X", x"0001", x"0002", x"000X", x"0010", x"0011", x"0012", x"001X", x"002", x"00X", x"0100", x"0101", x"0102", x"010X", x"011", x"012", x"01X", x"02", x"0X", x"1000", x"1001", x"1002", x"100X", x"101", x"102", x"10X", x"11", x"12", x"1X", x"2", x"X"),
		output_code => (16#0#, 16#37#, 16#1bf#, 16#6ff#, 16#1ffff#, 16#bf#, 16#4ff#, 16#ffff#, 16#1df#, 16#3df#, 16#7fff#, 16#27#, 16#3f#, 16#77f#, 16#27fff#, 16#fff#, 16#f#, 16#3bf#, 16#1ff#, 16#3ffff#, 16#2bf#, 16#2ff#, 16#2ffff#, 16#23f#, 16#13f#, 16#17fff#, 16#5f#, 16#25f#, 16#33fff#, 16#17#, 16#33f#, 16#ff#, 16#37fff#, 16#15f#, 16#67f#, 16#bfff#, 16#17ff#, 16#b#, 16#1b#, 16#35f#, 16#17f#, 16#2bfff#, 16#29f#, 16#7f#, 16#3fff#, 16#7ff#, 16#13#, 16#3b#, 16#df#, 16#57f#, 16#1bfff#, 16#19f#, 16#47f#, 16#23fff#, 16#21f#, 16#11f#, 16#1dfff#, 16#1bff#, 16#3#, 16#7#, 16#2df#, 16#37f#, 16#3bfff#, 16#39f#, 16#27f#, 16#13fff#, 16#31f#, 16#9f#, 16#3dfff#, 16#3ef#, 16#1f#, 16#dfff#, 16#bff#, 16#19#, 16#5#, 16#13ff#, 16#15#, 16#26f#, 16#16f#, 16#19fff#, 16#9#, 16#3ff#, 16#d#, 16#36f#, 16#ef#, 16#5fff#, 16#12f#, 16#3af#, 16#11fff#, 16#11#, 16#dff#, 16#1d#, 16#2ef#, 16#1ef#, 16#15fff#, 16#af#, 16#6f#, 16#9fff#, 16#2f#, 16#1af#, 16#1fff#, 16#1#, 16#5ff#),
		output_size => (1, 6, 10, 11, 18, 10, 11, 18, 10, 10, 18, 6, 10, 11, 18, 13, 6, 10, 11, 18, 10, 11, 18, 10, 10, 18, 10, 10, 18, 6, 10, 11, 18, 10, 11, 18, 13, 5, 6, 10, 11, 18, 10, 11, 18, 13, 5, 6, 10, 11, 18, 10, 11, 18, 10, 10, 18, 13, 5, 6, 10, 11, 18, 10, 11, 18, 10, 10, 18, 10, 10, 17, 13, 5, 5, 13, 5, 10, 10, 17, 5, 13, 5, 10, 10, 17, 9, 10, 17, 5, 12, 5, 10, 10, 17, 9, 10, 17, 9, 10, 17, 5, 12)
	);

	subtype hybrid_code_table11_t is hybrid_code_table_t (
		-- input_code(126 downto 0),
		output_code(126 downto 0),
		output_size(126 downto 0)
	);
	
	constant hybrid_code_table11_c : hybrid_code_table11_t := (
		-- input_code  => (x"0000000000000000", x"0000000000000001", x"0000000000000002", x"000000000000000X", x"000000000000001", x"000000000000002", x"00000000000000X", x"00000000000001", x"000000000000020", x"000000000000021", x"000000000000022", x"00000000000002X", x"0000000000000X", x"0000000000001", x"00000000000020", x"00000000000021", x"00000000000022", x"0000000000002X", x"000000000000X", x"000000000001", x"000000000002000", x"000000000002001", x"000000000002002", x"00000000000200X", x"00000000000201", x"00000000000202", x"0000000000020X", x"0000000000021", x"0000000000022", x"000000000002X", x"00000000000X", x"00000000001", x"00000000002", x"0000000000X", x"0000000001", x"0000000002", x"000000000X", x"000000001", x"000000002", x"00000000X", x"00000001", x"00000002", x"0000000X", x"00000010", x"00000011", x"00000012", x"0000001X", x"0000002", x"000000X", x"00000100", x"00000101", x"00000102", x"0000010X", x"0000011", x"0000012", x"000001X", x"000002", x"00000X", x"0000100", x"0000101", x"0000102", x"000010X", x"000011", x"000012", x"00001X", x"00002", x"0000X", x"0001000", x"0001001", x"0001002", x"000100X", x"000101", x"000102", x"00010X", x"00011", x"00012", x"0001X", x"0002", x"000X", x"0010000", x"0010001", x"0010002", x"001000X", x"001001", x"001002", x"00100X", x"00101", x"00102", x"0010X", x"0011", x"0012", x"001X", x"002", x"00X", x"01000000", x"01000001", x"01000002", x"0100000X", x"0100001", x"0100002", x"010000X", x"010001", x"010002", x"01000X", x"01001", x"01002", x"0100X", x"0101", x"0102", x"010X", x"011", x"012", x"01X", x"020", x"021", x"022", x"02X", x"0X", x"1", x"200", x"201", x"202", x"20X", x"21", x"22", x"2X", x"X"),
		output_code => (16#0#, 16#37#, 16#1f#, 16#3fff#, 16#17#, 16#4f#, 16#5fff#, 16#27#, 16#2f#, 16#9ff#, 16#5ff#, 16#7ffff#, 16#1fff#, 16#7#, 16#f#, 16#aff#, 16#6ff#, 16#3ffff#, 16#6fff#, 16#3b#, 16#6f#, 16#dff#, 16#3ff#, 16#fffff#, 16#eff#, 16#1ff#, 16#bffff#, 16#cff#, 16#2ff#, 16#dffff#, 16#2fff#, 16#2b#, 16#1b#, 16#4fff#, 16#33#, 16#b#, 16#fff#, 16#23#, 16#13#, 16#77ff#, 16#d#, 16#2d#, 16#37ff#, 16#1d#, 16#17f#, 16#57f#, 16#1ffff#, 16#5#, 16#17ff#, 16#3d#, 16#37f#, 16#77f#, 16#9ffff#, 16#2bf#, 16#6bf#, 16#cffff#, 16#39#, 16#27ff#, 16#25#, 16#1bf#, 16#5bf#, 16#2ffff#, 16#23f#, 16#63f#, 16#f7fff#, 16#19#, 16#7ff#, 16#15#, 16#3bf#, 16#7bf#, 16#affff#, 16#13f#, 16#53f#, 16#ffff#, 16#1df#, 16#5df#, 16#67fff#, 16#29#, 16#3bff#, 16#35#, 16#7f#, 16#47f#, 16#6ffff#, 16#33f#, 16#73f#, 16#8ffff#, 16#3df#, 16#7df#, 16#17fff#, 16#df#, 16#4df#, 16#47fff#, 16#11#, 16#1bff#, 16#3#, 16#ff#, 16#4ff#, 16#5ffff#, 16#27f#, 16#67f#, 16#effff#, 16#bf#, 16#4bf#, 16#4ffff#, 16#3f#, 16#43f#, 16#57fff#, 16#2df#, 16#6df#, 16#27fff#, 16#25f#, 16#65f#, 16#7fff#, 16#31#, 16#15f#, 16#55f#, 16#b7fff#, 16#2bff#, 16#1#, 16#9#, 16#35f#, 16#75f#, 16#77fff#, 16#5f#, 16#45f#, 16#37fff#, 16#bff#),
		output_size => (1, 6, 7, 15, 6, 7, 15, 6, 7, 12, 12, 20, 15, 6, 7, 12, 12, 20, 15, 6, 7, 12, 12, 20, 12, 12, 20, 12, 12, 20, 15, 6, 6, 15, 6, 6, 15, 6, 6, 15, 6, 6, 15, 6, 11, 11, 20, 6, 14, 6, 11, 11, 20, 11, 11, 20, 6, 14, 6, 11, 11, 20, 11, 11, 20, 6, 14, 6, 11, 11, 20, 11, 11, 20, 11, 11, 19, 6, 14, 6, 11, 11, 20, 11, 11, 20, 11, 11, 19, 11, 11, 19, 6, 14, 6, 11, 12, 20, 11, 11, 20, 11, 11, 20, 11, 11, 19, 11, 11, 19, 11, 11, 19, 6, 11, 11, 20, 14, 5, 6, 11, 11, 20, 11, 11, 20, 14)
	);

	subtype hybrid_code_table12_t is hybrid_code_table_t (
		-- input_code(108 downto 0),
		output_code(108 downto 0),
		output_size(108 downto 0)
	);
	
	constant hybrid_code_table12_c : hybrid_code_table12_t := (
		-- input_code  => (x"000000000000000000000000000", x"000000000000000000000000001", x"000000000000000000000000002", x"00000000000000000000000000X", x"00000000000000000000000001", x"00000000000000000000000002", x"0000000000000000000000000X", x"0000000000000000000000001", x"0000000000000000000000002", x"000000000000000000000000X", x"000000000000000000000001", x"000000000000000000000002", x"00000000000000000000000X", x"00000000000000000000001", x"00000000000000000000002", x"0000000000000000000000X", x"0000000000000000000001", x"0000000000000000000002", x"000000000000000000000X", x"000000000000000000001", x"000000000000000000002", x"00000000000000000000X", x"00000000000000000001", x"00000000000000000002", x"0000000000000000000X", x"0000000000000000001", x"0000000000000000002", x"000000000000000000X", x"000000000000000001", x"000000000000000002", x"00000000000000000X", x"00000000000000001", x"00000000000000002", x"0000000000000000X", x"0000000000000001", x"0000000000000002", x"000000000000000X", x"000000000000001", x"000000000000002", x"00000000000000X", x"00000000000001", x"00000000000002", x"0000000000000X", x"0000000000001", x"0000000000002", x"000000000000X", x"000000000001", x"000000000002", x"00000000000X", x"000000000010", x"000000000011", x"000000000012", x"00000000001X", x"00000000002", x"0000000000X", x"000000000100", x"000000000101", x"000000000102", x"00000000010X", x"00000000011", x"00000000012", x"0000000001X", x"0000000002", x"000000000X", x"000000001", x"000000002", x"00000000X", x"00000001", x"00000002", x"0000000X", x"0000001", x"0000002", x"000000X", x"000001", x"000002", x"00000X", x"00001", x"00002", x"0000X", x"0001", x"00020", x"00021", x"00022", x"0002X", x"000X", x"001", x"00200", x"00201", x"00202", x"0020X", x"0021", x"0022", x"002X", x"00X", x"01", x"02000", x"02001", x"02002", x"0200X", x"0201", x"0202", x"020X", x"021", x"022", x"02X", x"0X", x"1", x"2", x"X"),
		output_code => (16#0#, 16#3f#, 16#7f#, 16#ffff#, 16#1f#, 16#5f#, 16#7fff#, 16#2f#, 16#6f#, 16#bfff#, 16#f#, 16#4f#, 16#3fff#, 16#37#, 16#77#, 16#dfff#, 16#17#, 16#57#, 16#5fff#, 16#27#, 16#67#, 16#9fff#, 16#7#, 16#47#, 16#1fff#, 16#3b#, 16#7b#, 16#efff#, 16#1b#, 16#5b#, 16#6fff#, 16#2b#, 16#6b#, 16#afff#, 16#b#, 16#4b#, 16#2fff#, 16#33#, 16#73#, 16#cfff#, 16#13#, 16#53#, 16#4fff#, 16#23#, 16#63#, 16#fff#, 16#3d#, 16#7d#, 16#77ff#, 16#3#, 16#eff#, 16#13ff#, 16#bffff#, 16#5d#, 16#37ff#, 16#43#, 16#1ff#, 16#bff#, 16#7ffff#, 16#6ff#, 16#3ff#, 16#3ffff#, 16#1d#, 16#57ff#, 16#25#, 16#6d#, 16#17ff#, 16#5#, 16#2d#, 16#67ff#, 16#39#, 16#4d#, 16#27ff#, 16#19#, 16#d#, 16#47ff#, 16#29#, 16#15#, 16#7ff#, 16#9#, 16#55#, 16#cff#, 16#15ff#, 16#dffff#, 16#7bff#, 16#31#, 16#35#, 16#2ff#, 16#dff#, 16#fffff#, 16#8ff#, 16#19ff#, 16#9ffff#, 16#3bff#, 16#11#, 16#75#, 16#aff#, 16#1dff#, 16#1fffff#, 16#4ff#, 16#5ff#, 16#5ffff#, 16#ff#, 16#9ff#, 16#1ffff#, 16#5bff#, 16#1#, 16#21#, 16#1bff#),
		output_size => (1, 7, 8, 17, 7, 7, 16, 7, 7, 16, 7, 7, 16, 7, 7, 16, 7, 7, 16, 7, 7, 16, 7, 7, 16, 7, 7, 16, 7, 7, 16, 7, 7, 16, 7, 7, 16, 7, 7, 16, 7, 7, 16, 7, 7, 15, 7, 7, 15, 7, 12, 13, 20, 7, 15, 7, 12, 13, 20, 12, 13, 20, 7, 15, 6, 7, 15, 6, 7, 15, 6, 7, 15, 6, 7, 15, 6, 7, 15, 6, 7, 12, 13, 20, 15, 6, 7, 12, 13, 21, 12, 13, 20, 15, 6, 7, 12, 13, 21, 12, 13, 20, 12, 13, 20, 15, 6, 6, 15)
	);

	subtype hybrid_code_table13_t is hybrid_code_table_t (
		-- input_code(144 downto 0),
		output_code(144 downto 0),
		output_size(144 downto 0)
	);
	
	constant hybrid_code_table13_c : hybrid_code_table13_t := (
		-- input_code  => (x"0000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000001", x"00000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000001", x"0000000000000000000000000000000000000002", x"000000000000000000000000000000000000000X", x"000000000000000000000000000000000000001", x"000000000000000000000000000000000000002", x"00000000000000000000000000000000000000X", x"00000000000000000000000000000000000001", x"00000000000000000000000000000000000002", x"0000000000000000000000000000000000000X", x"0000000000000000000000000000000000001", x"0000000000000000000000000000000000002", x"000000000000000000000000000000000000X", x"000000000000000000000000000000000001", x"000000000000000000000000000000000002", x"00000000000000000000000000000000000X", x"00000000000000000000000000000000001", x"00000000000000000000000000000000002", x"0000000000000000000000000000000000X", x"0000000000000000000000000000000001", x"0000000000000000000000000000000002", x"000000000000000000000000000000000X", x"000000000000000000000000000000001", x"000000000000000000000000000000002", x"00000000000000000000000000000000X", x"00000000000000000000000000000001", x"00000000000000000000000000000002", x"0000000000000000000000000000000X", x"0000000000000000000000000000001", x"0000000000000000000000000000002", x"000000000000000000000000000000X", x"000000000000000000000000000001", x"000000000000000000000000000002", x"00000000000000000000000000000X", x"00000000000000000000000000001", x"00000000000000000000000000002", x"0000000000000000000000000000X", x"0000000000000000000000000001", x"0000000000000000000000000002", x"000000000000000000000000000X", x"000000000000000000000000001", x"000000000000000000000000002", x"00000000000000000000000000X", x"00000000000000000000000001", x"00000000000000000000000002", x"0000000000000000000000000X", x"0000000000000000000000001", x"0000000000000000000000002", x"000000000000000000000000X", x"000000000000000000000001", x"000000000000000000000002", x"00000000000000000000000X", x"00000000000000000000001", x"00000000000000000000002", x"0000000000000000000000X", x"0000000000000000000001", x"0000000000000000000002", x"000000000000000000000X", x"000000000000000000001", x"000000000000000000002", x"00000000000000000000X", x"00000000000000000001", x"00000000000000000002", x"0000000000000000000X", x"0000000000000000001", x"0000000000000000002", x"000000000000000000X", x"000000000000000001", x"000000000000000002", x"00000000000000000X", x"00000000000000001", x"00000000000000002", x"0000000000000000X", x"0000000000000001", x"0000000000000002", x"000000000000000X", x"000000000000001", x"000000000000002", x"00000000000000X", x"00000000000001", x"00000000000002", x"0000000000000X", x"0000000000001", x"0000000000002", x"000000000000X", x"000000000001", x"000000000002", x"00000000000X", x"00000000001", x"00000000002", x"0000000000X", x"0000000001", x"0000000002", x"000000000X", x"000000001", x"000000002", x"00000000X", x"00000001", x"00000002", x"0000000X", x"0000001", x"0000002", x"000000X", x"000001", x"000002", x"00000X", x"00001", x"00002", x"0000X", x"0001", x"0002", x"000X", x"001", x"002", x"00X", x"01", x"02", x"0X", x"100", x"101", x"102", x"10X", x"11", x"12", x"1X", x"2", x"X"),
		output_code => (16#0#, 16#7f#, 16#ff#, 16#ffff#, 16#3f#, 16#bf#, 16#7fff#, 16#5f#, 16#df#, 16#bfff#, 16#1f#, 16#9f#, 16#3fff#, 16#6f#, 16#ef#, 16#dfff#, 16#2f#, 16#af#, 16#5fff#, 16#4f#, 16#cf#, 16#9fff#, 16#f#, 16#8f#, 16#1fff#, 16#77#, 16#f7#, 16#efff#, 16#37#, 16#b7#, 16#6fff#, 16#57#, 16#d7#, 16#afff#, 16#17#, 16#97#, 16#2fff#, 16#67#, 16#e7#, 16#cfff#, 16#27#, 16#a7#, 16#4fff#, 16#47#, 16#c7#, 16#8fff#, 16#7#, 16#87#, 16#fff#, 16#7b#, 16#fb#, 16#f7ff#, 16#3b#, 16#bb#, 16#77ff#, 16#5b#, 16#db#, 16#b7ff#, 16#63#, 16#9b#, 16#37ff#, 16#23#, 16#1b#, 16#d7ff#, 16#43#, 16#eb#, 16#57ff#, 16#3#, 16#6b#, 16#97ff#, 16#7d#, 16#ab#, 16#17ff#, 16#3d#, 16#2b#, 16#e7ff#, 16#5d#, 16#cb#, 16#67ff#, 16#1d#, 16#4b#, 16#a7ff#, 16#6d#, 16#8b#, 16#27ff#, 16#2d#, 16#b#, 16#47ff#, 16#4d#, 16#f3#, 16#7ff#, 16#d#, 16#73#, 16#7bff#, 16#75#, 16#b3#, 16#3bff#, 16#35#, 16#33#, 16#5bff#, 16#55#, 16#d3#, 16#1bff#, 16#15#, 16#53#, 16#6bff#, 16#65#, 16#93#, 16#2bff#, 16#25#, 16#13#, 16#4bff#, 16#5#, 16#45#, 16#bff#, 16#39#, 16#79#, 16#73ff#, 16#19#, 16#59#, 16#33ff#, 16#29#, 16#69#, 16#53ff#, 16#9#, 16#49#, 16#13ff#, 16#31#, 16#71#, 16#63ff#, 16#61#, 16#11#, 16#23ff#, 16#41#, 16#21#, 16#43ff#, 16#51#, 16#5ff#, 16#dff#, 16#3ffff#, 16#1ff#, 16#9ff#, 16#1ffff#, 16#1#, 16#3ff#),
		output_size => (1, 8, 9, 17, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 7, 8, 16, 7, 8, 16, 7, 8, 16, 7, 8, 16, 7, 8, 16, 7, 8, 16, 7, 8, 16, 7, 8, 16, 7, 8, 16, 7, 8, 15, 7, 8, 15, 7, 8, 15, 7, 8, 15, 7, 8, 15, 7, 8, 15, 7, 8, 15, 7, 8, 15, 7, 8, 15, 7, 7, 15, 7, 7, 15, 7, 7, 15, 7, 7, 15, 7, 7, 15, 7, 7, 15, 7, 7, 15, 7, 7, 15, 7, 12, 12, 18, 12, 12, 18, 7, 15)
	);

	subtype hybrid_code_table14_t is hybrid_code_table_t (
		-- input_code(255 downto 0),
		output_code(255 downto 0),
		output_size(255 downto 0)
	);
	
	constant hybrid_code_table14_c : hybrid_code_table14_t := (
		-- input_code  => (x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000001", x"00000000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000001", x"0000000000000000000000000000000000000000002", x"000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000001", x"000000000000000000000000000000000000000002", x"00000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000001", x"00000000000000000000000000000000000000002", x"0000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000001", x"0000000000000000000000000000000000000002", x"000000000000000000000000000000000000000X", x"000000000000000000000000000000000000001", x"000000000000000000000000000000000000002", x"00000000000000000000000000000000000000X", x"00000000000000000000000000000000000001", x"00000000000000000000000000000000000002", x"0000000000000000000000000000000000000X", x"0000000000000000000000000000000000001", x"0000000000000000000000000000000000002", x"000000000000000000000000000000000000X", x"000000000000000000000000000000000001", x"000000000000000000000000000000000002", x"00000000000000000000000000000000000X", x"00000000000000000000000000000000001", x"00000000000000000000000000000000002", x"0000000000000000000000000000000000X", x"0000000000000000000000000000000001", x"0000000000000000000000000000000002", x"000000000000000000000000000000000X", x"000000000000000000000000000000001", x"000000000000000000000000000000002", x"00000000000000000000000000000000X", x"00000000000000000000000000000001", x"00000000000000000000000000000002", x"0000000000000000000000000000000X", x"0000000000000000000000000000001", x"0000000000000000000000000000002", x"000000000000000000000000000000X", x"000000000000000000000000000001", x"000000000000000000000000000002", x"00000000000000000000000000000X", x"00000000000000000000000000001", x"00000000000000000000000000002", x"0000000000000000000000000000X", x"0000000000000000000000000001", x"0000000000000000000000000002", x"000000000000000000000000000X", x"000000000000000000000000001", x"000000000000000000000000002", x"00000000000000000000000000X", x"00000000000000000000000001", x"00000000000000000000000002", x"0000000000000000000000000X", x"0000000000000000000000001", x"0000000000000000000000002", x"000000000000000000000000X", x"000000000000000000000001", x"000000000000000000000002", x"00000000000000000000000X", x"00000000000000000000001", x"00000000000000000000002", x"0000000000000000000000X", x"0000000000000000000001", x"0000000000000000000002", x"000000000000000000000X", x"000000000000000000001", x"000000000000000000002", x"00000000000000000000X", x"00000000000000000001", x"00000000000000000002", x"0000000000000000000X", x"0000000000000000001", x"0000000000000000002", x"000000000000000000X", x"000000000000000001", x"000000000000000002", x"00000000000000000X", x"00000000000000001", x"00000000000000002", x"0000000000000000X", x"0000000000000001", x"0000000000000002", x"000000000000000X", x"000000000000001", x"000000000000002", x"00000000000000X", x"00000000000001", x"00000000000002", x"0000000000000X", x"0000000000001", x"0000000000002", x"000000000000X", x"000000000001", x"000000000002", x"00000000000X", x"00000000001", x"00000000002", x"0000000000X", x"0000000001", x"0000000002", x"000000000X", x"000000001", x"000000002", x"00000000X", x"00000001", x"00000002", x"0000000X", x"0000001", x"0000002", x"000000X", x"000001", x"000002", x"00000X", x"00001", x"00002", x"0000X", x"0001", x"0002", x"000X", x"001", x"002", x"00X", x"01", x"02", x"0X", x"1", x"2", x"X"),
		output_code => (16#0#, 16#ff#, 16#1ff#, 16#1ffff#, 16#7f#, 16#17f#, 16#ffff#, 16#bf#, 16#1bf#, 16#17fff#, 16#3f#, 16#13f#, 16#7fff#, 16#df#, 16#1df#, 16#1bfff#, 16#5f#, 16#15f#, 16#bfff#, 16#9f#, 16#19f#, 16#13fff#, 16#1f#, 16#11f#, 16#3fff#, 16#ef#, 16#1ef#, 16#1dfff#, 16#6f#, 16#16f#, 16#dfff#, 16#af#, 16#1af#, 16#15fff#, 16#2f#, 16#12f#, 16#5fff#, 16#cf#, 16#1cf#, 16#19fff#, 16#4f#, 16#14f#, 16#9fff#, 16#8f#, 16#18f#, 16#11fff#, 16#f#, 16#10f#, 16#1fff#, 16#f7#, 16#1f7#, 16#1efff#, 16#77#, 16#177#, 16#efff#, 16#b7#, 16#1b7#, 16#16fff#, 16#37#, 16#137#, 16#6fff#, 16#ab#, 16#1d7#, 16#1afff#, 16#2b#, 16#d7#, 16#afff#, 16#cb#, 16#157#, 16#12fff#, 16#4b#, 16#57#, 16#2fff#, 16#8b#, 16#197#, 16#1cfff#, 16#b#, 16#97#, 16#cfff#, 16#f3#, 16#117#, 16#14fff#, 16#73#, 16#17#, 16#4fff#, 16#b3#, 16#1e7#, 16#18fff#, 16#33#, 16#e7#, 16#8fff#, 16#d3#, 16#167#, 16#10fff#, 16#53#, 16#67#, 16#fff#, 16#93#, 16#1a7#, 16#1f7ff#, 16#13#, 16#a7#, 16#f7ff#, 16#e3#, 16#127#, 16#177ff#, 16#63#, 16#27#, 16#77ff#, 16#a3#, 16#1c7#, 16#1b7ff#, 16#23#, 16#c7#, 16#b7ff#, 16#c3#, 16#147#, 16#137ff#, 16#43#, 16#47#, 16#37ff#, 16#83#, 16#187#, 16#1d7ff#, 16#3#, 16#87#, 16#d7ff#, 16#fd#, 16#107#, 16#57ff#, 16#7d#, 16#7#, 16#97ff#, 16#bd#, 16#1fb#, 16#17ff#, 16#3d#, 16#fb#, 16#e7ff#, 16#dd#, 16#17b#, 16#67ff#, 16#5d#, 16#7b#, 16#a7ff#, 16#9d#, 16#1bb#, 16#27ff#, 16#1d#, 16#bb#, 16#c7ff#, 16#ed#, 16#13b#, 16#47ff#, 16#6d#, 16#3b#, 16#87ff#, 16#ad#, 16#1db#, 16#7ff#, 16#2d#, 16#db#, 16#fbff#, 16#cd#, 16#15b#, 16#7bff#, 16#4d#, 16#5b#, 16#bbff#, 16#8d#, 16#19b#, 16#3bff#, 16#d#, 16#9b#, 16#dbff#, 16#f5#, 16#11b#, 16#5bff#, 16#75#, 16#1b#, 16#9bff#, 16#b5#, 16#1eb#, 16#1bff#, 16#35#, 16#eb#, 16#ebff#, 16#d5#, 16#16b#, 16#6bff#, 16#55#, 16#6b#, 16#abff#, 16#15#, 16#95#, 16#2bff#, 16#65#, 16#e5#, 16#cbff#, 16#25#, 16#a5#, 16#4bff#, 16#45#, 16#c5#, 16#8bff#, 16#5#, 16#85#, 16#bff#, 16#79#, 16#f9#, 16#f3ff#, 16#39#, 16#b9#, 16#73ff#, 16#59#, 16#d9#, 16#b3ff#, 16#19#, 16#99#, 16#33ff#, 16#69#, 16#e9#, 16#d3ff#, 16#29#, 16#a9#, 16#53ff#, 16#49#, 16#c9#, 16#93ff#, 16#9#, 16#89#, 16#13ff#, 16#71#, 16#f1#, 16#e3ff#, 16#31#, 16#b1#, 16#63ff#, 16#51#, 16#d1#, 16#a3ff#, 16#11#, 16#91#, 16#23ff#, 16#61#, 16#e1#, 16#c3ff#, 16#21#, 16#a1#, 16#43ff#, 16#41#, 16#c1#, 16#83ff#, 16#1#, 16#81#, 16#3ff#),
		output_size => (1, 9, 10, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 9, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 17, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 9, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16, 8, 8, 16)
	);

	subtype hybrid_code_table15_t is hybrid_code_table_t (
		-- input_code(256 downto 0),
		output_code(256 downto 0),
		output_size(256 downto 0)
	);
	
	constant hybrid_code_table15_c : hybrid_code_table15_t := (
		-- input_code  => (x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000000X", x"0000000000000000000000000000000000000000X", x"000000000000000000000000000000000000000X", x"00000000000000000000000000000000000000X", x"0000000000000000000000000000000000000X", x"000000000000000000000000000000000000X", x"00000000000000000000000000000000000X", x"0000000000000000000000000000000000X", x"000000000000000000000000000000000X", x"00000000000000000000000000000000X", x"0000000000000000000000000000000X", x"000000000000000000000000000000X", x"00000000000000000000000000000X", x"0000000000000000000000000000X", x"000000000000000000000000000X", x"00000000000000000000000000X", x"0000000000000000000000000X", x"000000000000000000000000X", x"00000000000000000000000X", x"0000000000000000000000X", x"000000000000000000000X", x"00000000000000000000X", x"0000000000000000000X", x"000000000000000000X", x"00000000000000000X", x"0000000000000000X", x"000000000000000X", x"00000000000000X", x"0000000000000X", x"000000000000X", x"00000000000X", x"0000000000X", x"000000000X", x"00000000X", x"0000000X", x"000000X", x"00000X", x"0000X", x"000X", x"00X", x"0X", x"X"),
		output_code => (16#0#, 16#1ff#, 16#ff#, 16#17f#, 16#7f#, 16#1bf#, 16#bf#, 16#13f#, 16#3f#, 16#1df#, 16#df#, 16#15f#, 16#5f#, 16#19f#, 16#9f#, 16#11f#, 16#1f#, 16#1ef#, 16#ef#, 16#16f#, 16#6f#, 16#1af#, 16#af#, 16#12f#, 16#2f#, 16#1cf#, 16#cf#, 16#14f#, 16#4f#, 16#18f#, 16#8f#, 16#10f#, 16#f#, 16#1f7#, 16#f7#, 16#177#, 16#77#, 16#1b7#, 16#b7#, 16#137#, 16#37#, 16#1d7#, 16#d7#, 16#157#, 16#57#, 16#197#, 16#97#, 16#117#, 16#17#, 16#1e7#, 16#e7#, 16#167#, 16#67#, 16#1a7#, 16#a7#, 16#127#, 16#27#, 16#1c7#, 16#c7#, 16#147#, 16#47#, 16#187#, 16#87#, 16#107#, 16#7#, 16#1fb#, 16#fb#, 16#17b#, 16#7b#, 16#1bb#, 16#bb#, 16#13b#, 16#3b#, 16#1db#, 16#db#, 16#15b#, 16#5b#, 16#19b#, 16#9b#, 16#11b#, 16#1b#, 16#1eb#, 16#eb#, 16#16b#, 16#6b#, 16#1ab#, 16#ab#, 16#12b#, 16#2b#, 16#1cb#, 16#cb#, 16#14b#, 16#4b#, 16#18b#, 16#8b#, 16#10b#, 16#b#, 16#1f3#, 16#f3#, 16#173#, 16#73#, 16#1b3#, 16#b3#, 16#133#, 16#33#, 16#1d3#, 16#d3#, 16#153#, 16#53#, 16#193#, 16#93#, 16#113#, 16#13#, 16#1e3#, 16#e3#, 16#163#, 16#63#, 16#1a3#, 16#a3#, 16#123#, 16#23#, 16#1c3#, 16#c3#, 16#143#, 16#43#, 16#183#, 16#83#, 16#103#, 16#3#, 16#1fd#, 16#fd#, 16#17d#, 16#7d#, 16#1bd#, 16#bd#, 16#13d#, 16#3d#, 16#1dd#, 16#dd#, 16#15d#, 16#5d#, 16#19d#, 16#9d#, 16#11d#, 16#1d#, 16#1ed#, 16#ed#, 16#16d#, 16#6d#, 16#1ad#, 16#ad#, 16#12d#, 16#2d#, 16#1cd#, 16#cd#, 16#14d#, 16#4d#, 16#18d#, 16#8d#, 16#10d#, 16#d#, 16#1f5#, 16#f5#, 16#175#, 16#75#, 16#1b5#, 16#b5#, 16#135#, 16#35#, 16#1d5#, 16#d5#, 16#155#, 16#55#, 16#195#, 16#95#, 16#115#, 16#15#, 16#1e5#, 16#e5#, 16#165#, 16#65#, 16#1a5#, 16#a5#, 16#125#, 16#25#, 16#1c5#, 16#c5#, 16#145#, 16#45#, 16#185#, 16#85#, 16#105#, 16#5#, 16#1f9#, 16#f9#, 16#179#, 16#79#, 16#1b9#, 16#b9#, 16#139#, 16#39#, 16#1d9#, 16#d9#, 16#159#, 16#59#, 16#199#, 16#99#, 16#119#, 16#19#, 16#1e9#, 16#e9#, 16#169#, 16#69#, 16#1a9#, 16#a9#, 16#129#, 16#29#, 16#1c9#, 16#c9#, 16#149#, 16#49#, 16#189#, 16#89#, 16#109#, 16#9#, 16#1f1#, 16#f1#, 16#171#, 16#71#, 16#1b1#, 16#b1#, 16#131#, 16#31#, 16#1d1#, 16#d1#, 16#151#, 16#51#, 16#191#, 16#91#, 16#111#, 16#11#, 16#1e1#, 16#e1#, 16#161#, 16#61#, 16#1a1#, 16#a1#, 16#121#, 16#21#, 16#1c1#, 16#c1#, 16#141#, 16#41#, 16#181#, 16#81#, 16#101#, 16#1#),
		output_size => (1, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9)
	);

end package hybrid_code_table;