library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.types_image.all;

-- Package Declaration Section
package hybrid_code_table is	

	type hybrid_flush_table_t is record
		-- active_prefix : array_unsigned_t;
		flush_word	: array_integer_t;
		flush_size	: array_integer_t;
	end record hybrid_flush_table_t;
	
	subtype hybrid_flush_table0_t is hybrid_flush_table_t (
		-- active_prefix(7 downto 0),
		flush_word(7 downto 0),
		flush_size(7 downto 0)
	);
	
	constant hybrid_flush_table0_c : hybrid_flush_table0_t := (
		-- active_prefix => (x"", x"0", x"01", x"02", x"4", x"44", x"7", x"8"),
		flush_word => (16#0#, 16#1#, 16#f#, 16#1f#, 16#3#, 16#3f#, 16#7#, 16#17#),
		flush_size => (1, 2, 5, 6, 3, 6, 5, 5)
	);

	subtype hybrid_flush_table1_t is hybrid_flush_table_t (
		-- active_prefix(12 downto 0),
		flush_word(12 downto 0),
		flush_size(12 downto 0)
	);
	
	constant hybrid_flush_table1_c : hybrid_flush_table1_t := (
		-- active_prefix => (x"", x"0", x"00", x"03", x"04", x"1", x"13", x"15", x"16", x"2", x"23", x"25", x"A"),
		flush_word => (16#0#, 16#1#, 16#7#, 16#17#, 16#37#, 16#5#, 16#f#, 16#5f#, 16#3f#, 16#3#, 16#2f#, 16#7f#, 16#1#),
		flush_size => (1, 3, 5, 6, 6, 3, 6, 7, 7, 3, 6, 7, 7)
	);

	subtype hybrid_flush_table2_t is hybrid_flush_table_t (
		-- active_prefix(12 downto 0),
		flush_word(12 downto 0),
		flush_size(12 downto 0)
	);
	
	constant hybrid_flush_table2_c : hybrid_flush_table2_t := (
		-- active_prefix => (x"", x"1", x"11", x"12", x"13", x"14", x"2", x"20", x"21", x"23", x"24", x"5", x"6"),
		flush_word => (16#0#, 16#1#, 16#b#, 16#1b#, 16#f#, 16#2f#, 16#5#, 16#7#, 16#17#, 16#1f#, 16#3f#, 16#3#, 16#13#),
		flush_size => (1, 3, 5, 5, 6, 6, 3, 5, 5, 6, 6, 5, 5)
	);

	subtype hybrid_flush_table3_t is hybrid_flush_table_t (
		-- active_prefix(16 downto 0),
		flush_word(16 downto 0),
		flush_size(16 downto 0)
	);
	
	constant hybrid_flush_table3_c : hybrid_flush_table3_t := (
		-- active_prefix => (x"", x"0", x"00", x"001", x"002", x"2", x"21", x"211", x"22", x"221", x"23", x"3", x"31", x"32", x"4", x"41", x"6"),
		flush_word => (16#0#, 16#1#, 16#b#, 16#5f#, 16#3f#, 16#5#, 16#17#, 16#7f#, 16#37#, 16#ff#, 16#4f#, 16#3#, 16#2f#, 16#6f#, 16#7#, 16#1f#, 16#f#),
		flush_size => (1, 3, 4, 7, 7, 3, 6, 8, 6, 8, 7, 4, 7, 7, 5, 7, 7)
	);

	subtype hybrid_flush_table4_t is hybrid_flush_table_t (
		-- active_prefix(12 downto 0),
		flush_word(12 downto 0),
		flush_size(12 downto 0)
	);
	
	constant hybrid_flush_table4_c : hybrid_flush_table4_t := (
		-- active_prefix => (x"", x"0", x"00", x"001", x"01", x"010", x"011", x"012", x"02", x"021", x"022", x"03", x"04"),
		flush_word => (16#0#, 16#1#, 16#3#, 16#37#, 16#b#, 16#f#, 16#2f#, 16#5f#, 16#7#, 16#3f#, 16#7f#, 16#17#, 16#1f#),
		flush_size => (1, 2, 4, 6, 4, 6, 6, 7, 5, 7, 7, 6, 7)
	);

	subtype hybrid_flush_table5_t is hybrid_flush_table_t (
		-- active_prefix(22 downto 0),
		flush_word(22 downto 0),
		flush_size(22 downto 0)
	);
	
	constant hybrid_flush_table5_c : hybrid_flush_table5_t := (
		-- active_prefix => (x"", x"2", x"20", x"200", x"2001", x"20010", x"2002", x"201", x"2010", x"20100", x"202", x"2020", x"21", x"210", x"2100", x"21000", x"211", x"212", x"22", x"220", x"2200", x"221", x"24"),
		flush_word => (16#0#, 16#1#, 16#5#, 16#b#, 16#4f#, 16#bf#, 16#2f#, 16#1b#, 16#6f#, 16#7f#, 16#3b#, 16#1f#, 16#3#, 16#7#, 16#17#, 16#ff#, 16#37#, 16#77#, 16#13#, 16#27#, 16#5f#, 16#f#, 16#3f#),
		flush_size => (1, 3, 3, 5, 7, 8, 7, 6, 7, 8, 6, 7, 5, 6, 6, 8, 7, 7, 5, 6, 7, 7, 8)
	);

	subtype hybrid_flush_table6_t is hybrid_flush_table_t (
		-- active_prefix(19 downto 0),
		flush_word(19 downto 0),
		flush_size(19 downto 0)
	);
	
	constant hybrid_flush_table6_c : hybrid_flush_table6_t := (
		-- active_prefix => (x"", x"0", x"00", x"000", x"0001", x"00010", x"0002", x"00020", x"001", x"0010", x"02", x"021", x"1", x"11", x"110", x"2", x"20", x"201", x"2010", x"3"),
		flush_word => (16#0#, 16#2#, 16#1#, 16#3#, 16#17#, 16#5f#, 16#37#, 16#3f#, 16#27#, 16#f#, 16#b#, 16#2f#, 16#5#, 16#7#, 16#6f#, 16#d#, 16#1b#, 16#1f#, 16#ff#, 16#7f#),
		flush_size => (2, 2, 3, 4, 6, 7, 6, 7, 6, 6, 5, 7, 4, 6, 7, 4, 5, 7, 8, 8)
	);

	subtype hybrid_flush_table7_t is hybrid_flush_table_t (
		-- active_prefix(15 downto 0),
		flush_word(15 downto 0),
		flush_size(15 downto 0)
	);
	
	constant hybrid_flush_table7_c : hybrid_flush_table7_t := (
		-- active_prefix => (x"", x"0", x"01", x"010", x"0101", x"0102", x"02", x"022", x"1", x"10", x"100", x"1001", x"1002", x"11", x"112", x"3"),
		flush_word => (16#0#, 16#1#, 16#b#, 16#17#, 16#df#, 16#3f#, 16#1b#, 16#5f#, 16#3#, 16#7#, 16#f#, 16#bf#, 16#7f#, 16#1f#, 16#1ff#, 16#ff#),
		flush_size => (1, 2, 5, 5, 8, 8, 5, 8, 4, 5, 5, 8, 8, 7, 9, 9)
	);

	subtype hybrid_flush_table8_t is hybrid_flush_table_t (
		-- active_prefix(28 downto 0),
		flush_word(28 downto 0),
		flush_size(28 downto 0)
	);
	
	constant hybrid_flush_table8_c : hybrid_flush_table8_t := (
		-- active_prefix => (x"", x"0", x"00", x"000", x"0000", x"00000", x"000000", x"0000000", x"00000000", x"000000000", x"0000000002", x"00000000020", x"00000001", x"000000010", x"00000002", x"0000002", x"00000020", x"00001", x"00002", x"0002", x"00020", x"00021", x"01", x"1", x"10", x"11", x"2", x"20", x"21"),
		flush_word => (16#0#, 16#2#, 16#6#, 16#1#, 16#5#, 16#d#, 16#3#, 16#13#, 16#b#, 16#1b#, 16#17f#, 16#ff#, 16#5f#, 16#bf#, 16#df#, 16#9f#, 16#3f#, 16#2f#, 16#1f#, 16#4f#, 16#6f#, 16#3ff#, 16#17#, 16#7#, 16#37#, 16#7f#, 16#27#, 16#f#, 16#1ff#),
		flush_size => (2, 3, 3, 3, 4, 4, 5, 5, 5, 5, 9, 9, 8, 8, 8, 8, 8, 7, 8, 7, 7, 10, 6, 6, 6, 9, 6, 7, 10)
	);

	subtype hybrid_flush_table9_t is hybrid_flush_table_t (
		-- active_prefix(33 downto 0),
		flush_word(33 downto 0),
		flush_size(33 downto 0)
	);
	
	constant hybrid_flush_table9_c : hybrid_flush_table9_t := (
		-- active_prefix => (x"", x"0", x"00", x"000", x"0000", x"00000", x"000000", x"0000000", x"00000000", x"000000000", x"0000000000", x"001", x"0001", x"00001", x"000000001", x"0000000001", x"00000000001", x"02", x"002", x"0000002", x"00000002", x"000000002", x"0010", x"00010", x"0000000010", x"00000000010", x"020", x"0020", x"00000020", x"000000020", x"00100", x"00000000100", x"0200", x"000000200"),
		flush_word => (16#0#, 16#1#, 16#2#, 16#3#, 16#8#, 16#9#, 16#a#, 16#b#, 16#c#, 16#1a#, 16#1b#, 16#47#, 16#74#, 16#76#, 16#1f#, 16#3f#, 16#ff#, 16#70#, 16#72#, 16#f5#, 16#f6#, 16#9f#, 16#75#, 16#77#, 16#bf#, 16#1ff#, 16#67#, 16#cf#, 16#ef#, 16#5f#, 16#f#, 16#7f#, 16#2f#, 16#df#),
		flush_size => (3, 3, 3, 3, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 8, 8, 9, 7, 7, 8, 8, 8, 7, 7, 8, 9, 7, 8, 8, 8, 7, 8, 8, 8)
	);

	subtype hybrid_flush_table10_t is hybrid_flush_table_t (
		-- active_prefix(33 downto 0),
		flush_word(33 downto 0),
		flush_size(33 downto 0)
	);
	
	constant hybrid_flush_table10_c : hybrid_flush_table10_t := (
		-- active_prefix => (x"", x"0", x"00", x"000", x"0000", x"00000", x"000000", x"0000000", x"00000000", x"1", x"01", x"001", x"00000001", x"000000001", x"00002", x"000002", x"0000002", x"00000002", x"000000002", x"10", x"010", x"000000010", x"0000000010", x"000020", x"0000020", x"00000020", x"000000020", x"100", x"0000000100", x"00000000100", x"0000200", x"00000200", x"00000001000", x"00002000"),
		flush_word => (16#0#, 16#1#, 16#2#, 16#3#, 16#4#, 16#5#, 16#c#, 16#d#, 16#e#, 16#f#, 16#f1#, 16#f3#, 16#19f#, 16#3f#, 16#6f#, 16#1ee#, 16#1f0#, 16#5f#, 16#13f#, 16#f2#, 16#f4#, 16#1fa#, 16#1fc#, 16#1ef#, 16#1f1#, 16#15f#, 16#1bf#, 16#af#, 16#1fd#, 16#1fe#, 16#9f#, 16#df#, 16#1ff#, 16#1df#),
		flush_size => (3, 3, 3, 3, 3, 3, 4, 4, 4, 8, 8, 8, 9, 9, 8, 9, 9, 9, 9, 8, 8, 9, 9, 9, 9, 9, 9, 8, 9, 9, 9, 9, 9, 9)
	);

	subtype hybrid_flush_table11_t is hybrid_flush_table_t (
		-- active_prefix(41 downto 0),
		flush_word(41 downto 0),
		flush_size(41 downto 0)
	);
	
	constant hybrid_flush_table11_c : hybrid_flush_table11_t := (
		-- active_prefix => (x"", x"0", x"00", x"000", x"0000", x"00000", x"000000", x"0000000", x"00000000", x"000000000", x"0000000000", x"00000000000", x"000000000000", x"0000000000000", x"00000000000000", x"000000000000000", x"01", x"001", x"0001", x"00001", x"000001", x"0000001", x"2", x"02", x"000000000002", x"0000000000002", x"00000000000002", x"010", x"0010", x"00010", x"000010", x"0000010", x"20", x"0000000000020", x"0100", x"00100", x"000100", x"00000000000200", x"01000", x"001000", x"010000", x"0100000"),
		flush_word => (16#0#, 16#1#, 16#2#, 16#3#, 16#4#, 16#5#, 16#6#, 16#7#, 16#8#, 16#9#, 16#a#, 16#b#, 16#c#, 16#d#, 16#e#, 16#f#, 16#1f#, 16#1f1#, 16#1f3#, 16#3df#, 16#33f#, 16#7f#, 16#3ec#, 16#3ed#, 16#37f#, 16#3fc#, 16#3fe#, 16#1f2#, 16#1f4#, 16#3f#, 16#bf#, 16#27f#, 16#1df#, 16#2ff#, 16#15f#, 16#23f#, 16#2bf#, 16#3ff#, 16#13f#, 16#1bf#, 16#3bf#, 16#17f#),
		flush_size => (4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 9, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 9, 9, 10, 10, 10, 10, 10, 9, 10, 10, 10, 10, 10, 10, 10)
	);

	subtype hybrid_flush_table12_t is hybrid_flush_table_t (
		-- active_prefix(35 downto 0),
		flush_word(35 downto 0),
		flush_size(35 downto 0)
	);
	
	constant hybrid_flush_table12_c : hybrid_flush_table12_t := (
		-- active_prefix => (x"", x"0", x"00", x"000", x"0000", x"00000", x"000000", x"0000000", x"00000000", x"000000000", x"0000000000", x"00000000000", x"000000000000", x"0000000000000", x"00000000000000", x"000000000000000", x"0000000000000000", x"00000000000000000", x"000000000000000000", x"0000000000000000000", x"00000000000000000000", x"000000000000000000000", x"0000000000000000000000", x"00000000000000000000000", x"000000000000000000000000", x"0000000000000000000000000", x"00000000000000000000000000", x"0000000001", x"00000000001", x"02", x"002", x"0002", x"00000000010", x"020", x"0020", x"0200"),
		flush_word => (16#0#, 16#1#, 16#2#, 16#3#, 16#4#, 16#a#, 16#b#, 16#c#, 16#d#, 16#e#, 16#f#, 16#10#, 16#11#, 16#12#, 16#13#, 16#14#, 16#15#, 16#16#, 16#17#, 16#18#, 16#19#, 16#1a#, 16#1b#, 16#1c#, 16#1d#, 16#1e#, 16#1f#, 16#1fc#, 16#1fd#, 16#1f8#, 16#1f9#, 16#1ff#, 16#ff#, 16#bf#, 16#3ff#, 16#1bf#),
		flush_size => (4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 6, 9, 9, 9, 9, 10, 9, 9, 10, 9)
	);

	subtype hybrid_flush_table13_t is hybrid_flush_table_t (
		-- active_prefix(47 downto 0),
		flush_word(47 downto 0),
		flush_size(47 downto 0)
	);
	
	constant hybrid_flush_table13_c : hybrid_flush_table13_t := (
		-- active_prefix => (x"", x"0", x"00", x"000", x"0000", x"00000", x"000000", x"0000000", x"00000000", x"000000000", x"0000000000", x"00000000000", x"000000000000", x"0000000000000", x"00000000000000", x"000000000000000", x"0000000000000000", x"00000000000000000", x"000000000000000000", x"0000000000000000000", x"00000000000000000000", x"000000000000000000000", x"0000000000000000000000", x"00000000000000000000000", x"000000000000000000000000", x"0000000000000000000000000", x"00000000000000000000000000", x"000000000000000000000000000", x"0000000000000000000000000000", x"00000000000000000000000000000", x"000000000000000000000000000000", x"0000000000000000000000000000000", x"00000000000000000000000000000000", x"000000000000000000000000000000000", x"0000000000000000000000000000000000", x"00000000000000000000000000000000000", x"000000000000000000000000000000000000", x"0000000000000000000000000000000000000", x"00000000000000000000000000000000000000", x"000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000", x"1", x"10"),
		flush_word => (16#0#, 16#1#, 16#2#, 16#3#, 16#4#, 16#5#, 16#6#, 16#7#, 16#8#, 16#9#, 16#a#, 16#b#, 16#c#, 16#d#, 16#e#, 16#f#, 16#10#, 16#11#, 16#24#, 16#25#, 16#26#, 16#27#, 16#28#, 16#29#, 16#2a#, 16#2b#, 16#2c#, 16#2d#, 16#2e#, 16#2f#, 16#30#, 16#31#, 16#32#, 16#33#, 16#34#, 16#35#, 16#36#, 16#37#, 16#38#, 16#39#, 16#3a#, 16#3b#, 16#3c#, 16#3d#, 16#3e#, 16#3f#, 16#7f#, 16#ff#),
		flush_size => (5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 8, 8)
	);

	subtype hybrid_flush_table14_t is hybrid_flush_table_t (
		-- active_prefix(84 downto 0),
		flush_word(84 downto 0),
		flush_size(84 downto 0)
	);
	
	constant hybrid_flush_table14_c : hybrid_flush_table14_t := (
		-- active_prefix => (x"", x"0", x"00", x"000", x"0000", x"00000", x"000000", x"0000000", x"00000000", x"000000000", x"0000000000", x"00000000000", x"000000000000", x"0000000000000", x"00000000000000", x"000000000000000", x"0000000000000000", x"00000000000000000", x"000000000000000000", x"0000000000000000000", x"00000000000000000000", x"000000000000000000000", x"0000000000000000000000", x"00000000000000000000000", x"000000000000000000000000", x"0000000000000000000000000", x"00000000000000000000000000", x"000000000000000000000000000", x"0000000000000000000000000000", x"00000000000000000000000000000", x"000000000000000000000000000000", x"0000000000000000000000000000000", x"00000000000000000000000000000000", x"000000000000000000000000000000000", x"0000000000000000000000000000000000", x"00000000000000000000000000000000000", x"000000000000000000000000000000000000", x"0000000000000000000000000000000000000", x"00000000000000000000000000000000000000", x"000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
		flush_word => (16#0#, 16#1#, 16#2#, 16#3#, 16#4#, 16#5#, 16#6#, 16#7#, 16#8#, 16#9#, 16#a#, 16#b#, 16#c#, 16#d#, 16#e#, 16#f#, 16#10#, 16#11#, 16#12#, 16#13#, 16#14#, 16#15#, 16#16#, 16#17#, 16#18#, 16#19#, 16#1a#, 16#1b#, 16#1c#, 16#1d#, 16#1e#, 16#1f#, 16#20#, 16#21#, 16#22#, 16#23#, 16#24#, 16#25#, 16#26#, 16#27#, 16#28#, 16#29#, 16#2a#, 16#56#, 16#57#, 16#58#, 16#59#, 16#5a#, 16#5b#, 16#5c#, 16#5d#, 16#5e#, 16#5f#, 16#60#, 16#61#, 16#62#, 16#63#, 16#64#, 16#65#, 16#66#, 16#67#, 16#68#, 16#69#, 16#6a#, 16#6b#, 16#6c#, 16#6d#, 16#6e#, 16#6f#, 16#70#, 16#71#, 16#72#, 16#73#, 16#74#, 16#75#, 16#76#, 16#77#, 16#78#, 16#79#, 16#7a#, 16#7b#, 16#7c#, 16#7d#, 16#7e#, 16#7f#),
		flush_size => (6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7)
	);

	subtype hybrid_flush_table15_t is hybrid_flush_table_t (
		-- active_prefix(255 downto 0),
		flush_word(255 downto 0),
		flush_size(255 downto 0)
	);
	
	constant hybrid_flush_table15_c : hybrid_flush_table15_t := (
		-- active_prefix => (x"", x"0", x"00", x"000", x"0000", x"00000", x"000000", x"0000000", x"00000000", x"000000000", x"0000000000", x"00000000000", x"000000000000", x"0000000000000", x"00000000000000", x"000000000000000", x"0000000000000000", x"00000000000000000", x"000000000000000000", x"0000000000000000000", x"00000000000000000000", x"000000000000000000000", x"0000000000000000000000", x"00000000000000000000000", x"000000000000000000000000", x"0000000000000000000000000", x"00000000000000000000000000", x"000000000000000000000000000", x"0000000000000000000000000000", x"00000000000000000000000000000", x"000000000000000000000000000000", x"0000000000000000000000000000000", x"00000000000000000000000000000000", x"000000000000000000000000000000000", x"0000000000000000000000000000000000", x"00000000000000000000000000000000000", x"000000000000000000000000000000000000", x"0000000000000000000000000000000000000", x"00000000000000000000000000000000000000", x"000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
		flush_word => (16#0#, 16#1#, 16#2#, 16#3#, 16#4#, 16#5#, 16#6#, 16#7#, 16#8#, 16#9#, 16#a#, 16#b#, 16#c#, 16#d#, 16#e#, 16#f#, 16#10#, 16#11#, 16#12#, 16#13#, 16#14#, 16#15#, 16#16#, 16#17#, 16#18#, 16#19#, 16#1a#, 16#1b#, 16#1c#, 16#1d#, 16#1e#, 16#1f#, 16#20#, 16#21#, 16#22#, 16#23#, 16#24#, 16#25#, 16#26#, 16#27#, 16#28#, 16#29#, 16#2a#, 16#2b#, 16#2c#, 16#2d#, 16#2e#, 16#2f#, 16#30#, 16#31#, 16#32#, 16#33#, 16#34#, 16#35#, 16#36#, 16#37#, 16#38#, 16#39#, 16#3a#, 16#3b#, 16#3c#, 16#3d#, 16#3e#, 16#3f#, 16#40#, 16#41#, 16#42#, 16#43#, 16#44#, 16#45#, 16#46#, 16#47#, 16#48#, 16#49#, 16#4a#, 16#4b#, 16#4c#, 16#4d#, 16#4e#, 16#4f#, 16#50#, 16#51#, 16#52#, 16#53#, 16#54#, 16#55#, 16#56#, 16#57#, 16#58#, 16#59#, 16#5a#, 16#5b#, 16#5c#, 16#5d#, 16#5e#, 16#5f#, 16#60#, 16#61#, 16#62#, 16#63#, 16#64#, 16#65#, 16#66#, 16#67#, 16#68#, 16#69#, 16#6a#, 16#6b#, 16#6c#, 16#6d#, 16#6e#, 16#6f#, 16#70#, 16#71#, 16#72#, 16#73#, 16#74#, 16#75#, 16#76#, 16#77#, 16#78#, 16#79#, 16#7a#, 16#7b#, 16#7c#, 16#7d#, 16#7e#, 16#7f#, 16#80#, 16#81#, 16#82#, 16#83#, 16#84#, 16#85#, 16#86#, 16#87#, 16#88#, 16#89#, 16#8a#, 16#8b#, 16#8c#, 16#8d#, 16#8e#, 16#8f#, 16#90#, 16#91#, 16#92#, 16#93#, 16#94#, 16#95#, 16#96#, 16#97#, 16#98#, 16#99#, 16#9a#, 16#9b#, 16#9c#, 16#9d#, 16#9e#, 16#9f#, 16#a0#, 16#a1#, 16#a2#, 16#a3#, 16#a4#, 16#a5#, 16#a6#, 16#a7#, 16#a8#, 16#a9#, 16#aa#, 16#ab#, 16#ac#, 16#ad#, 16#ae#, 16#af#, 16#b0#, 16#b1#, 16#b2#, 16#b3#, 16#b4#, 16#b5#, 16#b6#, 16#b7#, 16#b8#, 16#b9#, 16#ba#, 16#bb#, 16#bc#, 16#bd#, 16#be#, 16#bf#, 16#c0#, 16#c1#, 16#c2#, 16#c3#, 16#c4#, 16#c5#, 16#c6#, 16#c7#, 16#c8#, 16#c9#, 16#ca#, 16#cb#, 16#cc#, 16#cd#, 16#ce#, 16#cf#, 16#d0#, 16#d1#, 16#d2#, 16#d3#, 16#d4#, 16#d5#, 16#d6#, 16#d7#, 16#d8#, 16#d9#, 16#da#, 16#db#, 16#dc#, 16#dd#, 16#de#, 16#df#, 16#e0#, 16#e1#, 16#e2#, 16#e3#, 16#e4#, 16#e5#, 16#e6#, 16#e7#, 16#e8#, 16#e9#, 16#ea#, 16#eb#, 16#ec#, 16#ed#, 16#ee#, 16#ef#, 16#f0#, 16#f1#, 16#f2#, 16#f3#, 16#f4#, 16#f5#, 16#f6#, 16#f7#, 16#f8#, 16#f9#, 16#fa#, 16#fb#, 16#fc#, 16#fd#, 16#fe#, 16#ff#),
		flush_size => (8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8)
	);

end package hybrid_code_table;